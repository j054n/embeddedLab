`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:24:17 03/12/2014 
// Design Name: 
// Module Name:    lab4Control 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab4Control(
    input CLK,
    input dataAvailable,
    output loadFirstSign,
    output loadFirstDigit,
    output loadSecondDigit,
    output loadSecondSign,
    output addNumbers,
    output displayAnswer,
	 output dataReady
	 
    );


endmodule
