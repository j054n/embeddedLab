`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:28:04 03/12/2014 
// Design Name: 
// Module Name:    lab4DataPath 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab4DataPath(
    input [7:0] dataIn,
    output [7:0] dataOut,
    input loadFirstSign,
    input loadFirstDigit,
    input loadSecondDigit,
    input loadSecondSign,
    input addNumbers,
    input displayAnswer,
    input CLK
    );



endmodule
