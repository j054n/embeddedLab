`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:19:21 03/12/2014 
// Design Name: 
// Module Name:    asciiTo4BitBinary 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module asciiTo4BitBinary(
    input [7:0] input8BitAscii,
    output [3:0] output4BitBinary
    );


endmodule
