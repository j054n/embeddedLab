`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:22:24 03/12/2014 
// Design Name: 
// Module Name:    binary16BitTo4DigitHex 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module binary16BitTo4DigitHex(
    input [15:0] inputBinary16Bit,
    output hexDigit0,
    output hexDigit1,
    output hexDigit2,
    output hexDigit3
    );


endmodule
