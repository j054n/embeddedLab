//
// lab1 : version 08/29/2012
//                  
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
//////////////////////////////////////////////////////////////////////////////////
module gates(
    input A0,
    input B0,
    output F0,
    input A1,
    input B1,
    output F1,
    input A2,
    input B2,
    output F2,
    input A3,
    input B3,
    output F3
    );

	// Write code starting here ...

endmodule
