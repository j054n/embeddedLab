//
// lab2 : version 09/04/2012
//                  
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module op_4bit(
    input [3:0] d,
    output parity
    );

	// design parity as sum of products

endmodule
