`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module nextupcount3(
    input [2:0] q,
    output [2:0] next_q
    );

endmodule
