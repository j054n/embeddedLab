`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:06:34 03/13/2014 
// Design Name: 
// Module Name:    addTwoNumbers 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module addTwoNumbers(
    input [15:0] NumberA,
    input [15:0] NumberB,
    output [15:0] Result
    );


endmodule
